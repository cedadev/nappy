netcdf \4010 {
dimensions:
	time = 2 ;
	altitude = 2 ;
	latitude = 7 ;
	longitude = 13 ;
variables:
	double time(time) ;
		time:name = "time (hours since 1980-06-01 00:00:00)" ;
		time:long_name = "time (hours since 1980-06-01 00:00:00)" ;
		time:standard_name = "time" ;
		time:units = "hours since 1980-06-01 00:00:00" ;
		time:calendar = "gregorian" ;
		time:axis = "T" ;
	double altitude(altitude) ;
		altitude:units = "km" ;
		altitude:long_name = "Altitude (km)" ;
		altitude:name = "Altitude" ;
	double latitude(latitude) ;
		latitude:units = "degrees_north" ;
		latitude:long_name = "Latitude (degrees_north)" ;
		latitude:standard_name = "latitude" ;
		latitude:name = "Latitude" ;
		latitude:axis = "Y" ;
	double longitude(longitude) ;
		longitude:modulo = 360. ;
		longitude:name = "Longitude" ;
		longitude:long_name = "Latitude (degrees_east)" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:axis = "X" ;
		longitude:topology = "circular" ;
	double temperature(time, altitude, latitude, longitude) ;
		temperature:title = "Temperature" ;
		temperature:long_name = "Temperature" ;
		temperature:units = "K" ;
		temperature:missing_value = 1000. ;
		temperature:nasa_ames_var_number = 0 ;

// global attributes:
		:Conventions = "CF-1.0" ;
		:comment = "==== Special Comments follow ====\nExample of FFI 4010.\nThis example illustrating NASA Ames file format index 4010 is entirely fictitious.\nData have been made up for the purpose of illustrating the use of the format. They\nconsist in an imaginary calculated temperature distribution over a longitude-lati-\ntude-altitude grid at 6 o\'clock and noon on the 21st of June 1980. The grid is\ndefined in lines 8, 9, 11, 12 and 13. Longitude ranges from 30 degrees West to 30\ndegrees East by intervals of 5 degrees. Latitude ranges from 90 North to 90 South by\nnegative intervals of 30 degrees. Altitude takes the two values of 20 and 50 km.\nIf the temperature is written as T(lon, lat, alt, time), the record below thus reads,\nfor each of the two times t = 6 and t = 12,\nt\nT(-30, 90, 20, t) . . . T(30, 90, 20, t)\n. . .                   . . .\nT(-30, -90, 20, t). . . T(30, -90, 20, t)\nT(-30, 90, 50, t) . . . T(30, 90, 50, t)\n. . .                   . . .\nT(-30, -90, 50, t). . . T(30, -90, 50, t)\n==== Special Comments end ====\n==== Normal Comments follow ====\nThe files included in this data set illustrate each of the 9 NASA Ames file format\nindices (FFI). A detailed description of the NASA Ames format can be found on the Web\nsite of the British Atmospheric Data Centre (BADC) at\nhttp://www.badc.rl.ac.uk/help/formats/NASA-Ames/\nE-mail contact: badc@rl.ac.uk\nReference: S. E. Gaines and R. S. Hipskind, Format Specification for Data Exchange,\nVersion 1.3, 1998. This work can be found at\nhttp://cloud1.arc.nasa.gov/solve/archiv/archive.tutorial.html and a copy of it at\nhttp://www.badc.rl.ac.uk/help/formats/NASA-Ames/G-and-H-June-1998.html\n==== Normal Comments end ====" ;
		:title = "NERC Data Grid (NDG) project" ;
		:file_number_in_set = 13 ;
		:source = "Imaginary 3-D stratospheric radiative model" ;
		:first_valid_date_of_data = 1980, 6, 21 ;
		:total_files_in_set = 13 ;
		:no_of_nasa_ames_header_lines = 53 ;
		:file_format_index = 4010 ;
		:institution = "De Rudder, Anne (ONAME from NASA Ames file); Rutherford Appleton Laboratory, Chilton OX11 0QX, UK - Tel.: +44 (0) 1235 445837 (ORG from NASA Ames file)." ;
		:history = "2002-10-31 - NASA Ames File created/revised.\n\n2021-05-10 15:14:45 - Converted to CDMS (NetCDF) format using nappy-0.3.0." ;
data:

 time = 6, 12 ;

 altitude = 20, 50 ;

 latitude = 90, 60, 30, 0, -30, -60, -90 ;

 longitude = -30, -25, -20, -15, -10, -5, 0, 5, 10, 15, 20, 25, 30 ;

 temperature =
  230, 230, 230, 230, 230, 230, 230, 230, 230, 230, 230, 230, 230,
  216, 216.5, 217, 218, 218.5, 219, 220, 220.4, 220.4, 220.9, 221.3, 221, 
    220.7,
  210.6, 211, 211.4, 211.8, 212.2, 212.6, 213, 213, 213.1, 213, 213.5, 213, 
    213.1,
  205.4, 206, 206.6, 207.2, 207.8, 208.4, 209, 209.2, 209.8, 210.3, 210, 
    209.8, 209.7,
  204, 204.6, 205, 205.7, 206.2, 206.8, 207, 207.4, 207.8, 208.2, 208.6, 
    208.3, 208,
  194.7, 195.2, 196, 196.6, 197.2, 197.5, 198, 198.4, 198.7, 198.9, 199.3, 
    199.5, 199.1,
  185, 185, 185, 185, 185, 185, 185, 185, 185, 185, 185, 185, 185,
  260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260,
  230, 230.5, 231, 233, 233.7, 234.2, 235, 235.5, 236, 236.5, 237, 237.5, 238,
  217.6, 218.3, 219, 219.3, 219.7, 220, 225, 225.8, 226.4, 227, 227.8, 228.5, 
    229.1,
  216.2, 216.7, 217, 217.4, 218.1, 218.5, 219, 219.8, 221, 221.6, 222, 223, 
    224,
  212.1, 212.7, 213, 213.5, 213.7, 214, 214, 214.5, 215.1, 216, 217, 218, 219,
  198.4, 199, 199.4, 200, 200.6, 201.1, 201, 201.5, 202, 202.8, 203.4, 204, 
    205,
  183, 183, 183, 183, 183, 183, 183, 183, 183, 183, 183, 183, 183,
  240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240,
  228.6, 228.7, 228.8, 229, 229.3, 229.8, 230, 230.5, 231, 231.5, 232, 231.5, 
    231,
  221.3, 221.7, 222, 222.4, 222.6, 223, 223, 223.6, 224, 224.4, 225, 224.5, 
    224,
  216.8, 217, 217.3, 217.8, 218, 218.4, 219, 219.3, 219.6, 220.3, 220.8, 
    219.9, 219,
  215.1, 215.4, 215.7, 216, 216.3, 216.6, 217, 217.5, 218, 218.6, 219, 218.9, 
    218.4,
  207.4, 207.5, 207.6, 207.7, 207.8, 207.9, 208, 208.2, 208.4, 208.6, 208.3, 
    208, 208.3,
  195, 195, 195, 195, 195, 195, 195, 195, 195, 195, 195, 195, 195,
  270, 270, 270, 270, 270, 270, 270, 270, 270, 270, 270, 270, 270,
  243, 243.5, 244, 244.3, 244.7, 245, 245, 245.2, 245.5, 250, 250.8, 251, 251,
  232.1, 232.7, 233, 234, 234.3, 234.7, 235, 235.3, 235.7, 236.2, 236.8, 
    236.6, 236.1,
  226.4, 226.8, 227, 227.4, 228, 228.8, 229, 229.8, 229.7, 230.3, 230.4, 
    230.3, 230,
  222.7, 222.8, 222.9, 223.2, 223.5, 224, 224, 224.5, 225, 225.2, 225.3, 225, 
    224.9,
  209.8, 210, 210.2, 210.4, 210.6, 210.8, 211, 211, 211.2, 211.3, 212, 212.1, 
    211.8,
  193, 193, 193, 193, 193, 193, 193, 193, 193, 193, 193, 193, 193 ;
}
